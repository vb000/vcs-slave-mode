module hello;
  
  initial begin
    $display("Hello!\n");
  end

endmodule
